.title KiCad schematic
.include "C:/AE/MAX16832C/_models/B3100.spice.txt"
.include "C:/AE/MAX16832C/_models/C2012X7R2A104K125AA_p.mod"
.include "C:/AE/MAX16832C/_models/C2012X7R2E103K125AA_p.mod"
.include "C:/AE/MAX16832C/_models/C3216X7R2E104K160AA_p.mod"
.include "C:/AE/MAX16832C/_models/C3225X7R2A105K200AA_p.mod"
.include "C:/AE/MAX16832C/_models/MAX16832C.LIB"
.include "C:/AE/MAX16832C/_models/PD_1210_7447709221_220u.lib"
.include "C:/AE/MAX16832C/_models/XLamp-XML-spice.txt"
.include "C:/AE/MAX16832C/_models/ntc_20130313.lib"
V2 /CTRL 0 PULSE(0 {VPUL} {DELAY} {TR} {TF} {DUTY} {CYCLE})
XU1 /A VCC 0 0 /LX /CTRL /TEMP MAX16832C
XU4 VCC 0 C3225X7R2A105K200AA_p
XU2 VCC 0 C2012X7R2A104K125AA_p
XU7 /LX /K PD_1210_7447709221_220u
R2 VCC /A {RSNS}
D1 /LX VCC DI_B3100
R3 VCC /A {RSNS}
XU6 /A /K C3216X7R2E104K160AA_p
D2 /A /B1 XM
D3 /B1 /B2 XM
D4 /B2 /B3 XM
D5 /B3 /B4 XM
D6 /B4 /B5 XM
D7 /B5 /K XM
XU3 /NTC 0 C2012X7R2E103K125AA_p
XU5 /NTC 0 B57452V5104J062
V1 VCC 0 {VSOURCE}
R1 /TEMP /NTC {RNTC}
.end
